package pkg;

  //-----------------------------------------------------
  // Interfaces
  //-----------------------------------------------------
  //`include "mem_if.sv"


  //-----------------------------------------------------
  // cLasses
  //-----------------------------------------------------
  `include "transaction.sv"

  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "subscriber.sv"

  `include "env.sv"


endpackage