// classes (inside pkg.svh)
`include "transaction.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "subscriber.sv"
`include "env.sv"
// interfaces
`include "mem_if.sv"

//
module memory16_32_tb //import pkg::*;
  ();


  //================================================================//
  //======================    PARAMETERS    ========================//
  //================================================================//
  localparam clk_period = 4;


  //================================================================//
  //======================    PORTS DECLARTION    ==================//
  //================================================================//
  logic                     i_mem_clk;
  logic                     i_mem_rst_n;


  //================================================================//
  //======================    Interfaces  ==========================//
  //================================================================//
  mem_if dut_if(i_mem_clk, i_mem_rst_n);
  virtual mem_if vif;


  //================================================================//
  //======================    DUT  =================================//
  //================================================================//
  memory16_32 DUT ( 
      dut_if
    );


  //================================================================//
  //======================    Classes  =============================//
  //================================================================//
  env ENV;


  //================================================================//
  //======================    Tests    =============================//
  //================================================================//
  initial begin
    i_mem_clk   = 0;
    i_mem_rst_n = 0;
    
    // Reset
    repeat (2) @(posedge i_mem_clk) i_mem_rst_n = 0;
    i_mem_rst_n = 1;
    
    // Interface
    vif = dut_if;

    // Enviroment
    ENV = new(vif);
    ENV.build();
    ENV.run();

  end


  //================================================================//
  //======================    CLOCK    =============================//
  //================================================================//
  always #(clk_period*0.5) i_mem_clk = ~i_mem_clk;


  //================================================================//
  //================================================================//
  //================================================================//


endmodule
